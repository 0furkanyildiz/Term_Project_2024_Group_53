library verilog;
use verilog.vl_types.all;
entity SSCDM_vlg_vec_tst is
end SSCDM_vlg_vec_tst;
